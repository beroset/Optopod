.title KiCad schematic
.include "/home/ejb/spice_models/APTD3216P3C-P22.lib"
.include "/home/ejb/spice_models/APTD3216SF4C-P22.lib"
.include "/home/ejb/spice_models/BC817-40.lib"
VJ1 +3V3 GND dc 3.3
Vin1 TX1 GND pulse(0 3.3 0.1u 0.1u 0.1u 1u 2u)
XQ3 Net-_Q2-Pad1_ Net-_Q3-Pad1_ GND BC817-40
R3 Net-_Q3-Pad1_ TX1 5.1k
R2 +3V3 Net-_Q2-Pad1_ 330
R5 Net-_Q3-Pad1_ GND 1.5k
XQ4 +3V3 Net-_Q4-Pad1_ Net-_Q4-Pad2_ BC817-40
R9 Net-_Q4-Pad2_ Net-_D2-Pad2_ 91
D2 Net-_D2-Pad2_ GND APTD3216SF4C-P22
XQ6 Net-_Q4-Pad1_ Net-_Q6-Pad1_ GND BC817-40
R8 Net-_Q6-Pad1_ TX2 5.1k
R7 +3V3 Net-_Q4-Pad1_ 330
R10 Net-_Q6-Pad1_ GND 1.5k
D1 Net-_D1-Pad2_ GND APTD3216SF4C-P22
R4 Net-_Q2-Pad2_ Net-_D1-Pad2_ 91
XQ2 +3V3 Net-_Q2-Pad1_ Net-_Q2-Pad2_ BC817-40
.tran 1n 4u 
.end
